library verilog;
use verilog.vl_types.all;
entity lab4_individual_vlg_vec_tst is
end lab4_individual_vlg_vec_tst;
