library verilog;
use verilog.vl_types.all;
entity counter8_vlg_vec_tst is
end counter8_vlg_vec_tst;
