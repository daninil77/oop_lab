library verilog;
use verilog.vl_types.all;
entity d_latch_vlg_vec_tst is
end d_latch_vlg_vec_tst;
