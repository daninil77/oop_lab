library verilog;
use verilog.vl_types.all;
entity secundomer_vlg_vec_tst is
end secundomer_vlg_vec_tst;
