library verilog;
use verilog.vl_types.all;
entity synchronizer_vlg_vec_tst is
end synchronizer_vlg_vec_tst;
