library verilog;
use verilog.vl_types.all;
entity shift_reg_left_4_vlg_vec_tst is
end shift_reg_left_4_vlg_vec_tst;
