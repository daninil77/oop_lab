library verilog;
use verilog.vl_types.all;
entity dff_rse_vlg_vec_tst is
end dff_rse_vlg_vec_tst;
