library verilog;
use verilog.vl_types.all;
entity rs_trig_nand_vlg_vec_tst is
end rs_trig_nand_vlg_vec_tst;
